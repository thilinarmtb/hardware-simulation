`define DEFAULT_WIDTH 12
