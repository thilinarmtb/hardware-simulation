`define DEFAULT_WIDTH 8
